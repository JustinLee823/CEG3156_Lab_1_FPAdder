library verilog;
use verilog.vl_types.all;
entity sevenBitUpCounter_vlg_vec_tst is
end sevenBitUpCounter_vlg_vec_tst;
