library ieee;
use ieee.std_logic_1164.all;

entity tenBitAdder is
	port(i_a, i_b : in std_logic_vector(9 downto 0);
		i_cin : in std_logic;
		o_cout : out std_logic;
		o_overflow : out std_logic;
		o_Value : out std_logic_vector(8 downto 0));
end tenBitAdder;

architecture rtl of tenBitAdder is

	signal carry : std_logic_vector(10 downto 0);
	signal sign_a, sign_b : std_logic;
	
begin
	sign_a <= i_a(9);
	sign_b <= i_b(9);
	carry(0) <= i_cin;
	
	o_Value(0) <= i_a(0) xor i_b(0) xor carry(0);
	o_Value(1) <= i_a(1) xor i_b(1) xor carry(1);
	o_Value(2) <= i_a(2) xor i_b(2) xor carry(2);
	o_Value(3) <= i_a(3) xor i_b(3) xor carry(3);
	o_Value(4) <= i_a(4) xor i_b(4) xor carry(4);
	o_Value(5) <= i_a(5) xor i_b(5) xor carry(5);
	o_Value(6) <= i_a(6) xor i_b(6) xor carry(6);
	o_Value(7) <= i_a(7) xor i_b(7) xor carry(7);
	o_Value(8) <= i_a(8) xor i_b(8) xor carry(8);
	
	
	
	carry(1) <= (i_a(0) and i_b(0)) or (i_a(0) and carry(0)) or (i_b(0) and  carry(0));
	carry(2) <= (i_a(1) and i_b(1)) or (i_a(1) and carry(1)) or (i_b(1) and  carry(1));
	carry(3) <= (i_a(2) and i_b(2)) or (i_a(2) and carry(2)) or (i_b(2) and  carry(2));
	carry(4) <= (i_a(3) and i_b(3)) or (i_a(3) and carry(3)) or (i_b(3) and  carry(3));
	carry(5) <= (i_a(4) and i_b(4)) or (i_a(4) and carry(4)) or (i_b(4) and  carry(4));
	carry(6) <= (i_a(5) and i_b(5)) or (i_a(5) and carry(5)) or (i_b(5) and  carry(5));
	carry(7) <= (i_a(6) and i_b(6)) or (i_a(6) and carry(6)) or (i_b(6) and  carry(6));
	carry(8) <= (i_a(7) and i_b(7)) or (i_a(7) and carry(7)) or (i_b(7) and  carry(7));
	carry(9) <= (i_a(8) and i_b(8)) or (i_a(8) and carry(8)) or (i_b(8) and  carry(8));
	carry(10) <= (i_a(9) and i_b(9)) or (i_a(9) and carry(9)) or (i_b(9) and carry(9));
	
	o_overflow <= carry(10) xor carry(9);
	o_cout <= carry(10);
end rtl;