LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY eightBitShiftRegister IS
	PORT(
		i_resetBar, i_load	: IN	STD_LOGIC;
		i_clock			: IN	STD_LOGIC;
		i_Value			: IN	STD_LOGIC_VECTOR(7 downto 0);
		o_Value			: OUT	STD_LOGIC_VECTOR(7 downto 0));
END eightBitShiftRegister;

ARCHITECTURE rtl OF eightBitShiftRegister IS
	SIGNAL int_Value, int_notValue : STD_LOGIC_VECTOR(7 downto 0);

	COMPONENT enARdFF_2
		PORT(
			i_resetBar	: IN	STD_LOGIC;
			i_d		: IN	STD_LOGIC;
			i_enable	: IN	STD_LOGIC;
			i_clock		: IN	STD_LOGIC;
			o_q, o_qBar	: OUT	STD_LOGIC);
	END COMPONENT;

BEGIN

	dff7 : enARdFF_2
	port map(
		i_resetBar => i_resetBar,
		i_clock => i_clock,
		i_enable => i_load, 
		i_d => i_Value(0),
		o_q => int_Value(7),
		o_qBar => int_notValue(7));

	dff6 : enARdFF_2
	port map(
		i_resetBar => i_resetBar,
		i_clock => i_clock,
		i_enable => i_load, 
		i_d => i_Value(7),
		o_q => int_Value(6),
		o_qBar => int_notValue(6));

	dff5 : enARdFF_2
	port map(
		i_resetBar => i_resetBar,
		i_clock => i_clock,
		i_enable => i_load, 
		i_d => i_Value(6),
		o_q => int_Value(5),
		o_qBar => int_notValue(5));	

	dff4 : enARdFF_2
	port map(
		i_resetBar => i_resetBar,
		i_clock => i_clock,
		i_enable => i_load, 
		i_d => i_Value(5),
		o_q => int_Value(4),
		o_qBar => int_notValue(4));

	dff3 : enARdFF_2
	port map(
		i_resetBar => i_resetBar,
		i_clock => i_clock,
		i_enable => i_load, 
		i_d => i_Value(4),
		o_q => int_Value(3),
		o_qBar => int_notValue(3));

	dff2 : enARdFF_2
	port map(
		i_resetBar => i_resetBar,
		i_clock => i_clock,
		i_enable => i_load,
		i_d => i_Value(3),
		o_q => int_Value(2),
		o_qBar => int_notValue(2));

	dff1 : enARdFF_2
	port map(
		i_resetBar => i_resetBar,
		i_clock => i_clock,
		i_enable => i_load,
		i_d => i_Value(2),
		o_q => int_Value(1),
		o_qBar => int_notValue(1));	

	dff0 : enARdFF_2
	port map(
		i_resetBar => i_resetBar,
		i_clock => i_clock,
		i_enable => i_load,
		i_d => i_Value(1),
		o_q => int_Value(0),
		o_qBar => int_notValue(0));	
	
	o_Value <= int_Value;
END rtl;